module tab();
	initial begin
		$display("HH:%b", 8'b11111111);
		$display("SD:%b", 8'b00001000);
		$display("BD:%b", 8'b10001000);
	end
endmodule
