module tab();
	initial begin
		$display("HH:%b", 4'b11111111);
		$display("SD:%b", 4'b00001000);
		$display("BD:%b", 4'b10001000);
	end
endmodule
